module top(

    input logic Clk, 
    input logic Reset, 
    input logic Walk, 

    output logic [2:0] LED 

); 




// https://docs.google.com/document/d/1k-O6FEl9OJP1CAzrinxhXka3euEQgAkbo8tkSL4IqJI/edit


endmodule 
